module incrementor
(
	input 		[63:0]	a		,
	output 		[63:0]	b
);
	
	assign 		b 		= a+1;

endmodule
